library ieee;
use ieee.std_logic_1164.all;
entity gaire_reduced_xor is
	port(
	a: in std_logic_vector(7 downto 0);
	y: out std_logic);
end gaire_reduced_xor;

architecture cascade1_arch of gaire_reduced_xor is
begin
	y <= a(0) xor a(1) xor a(2) xor a(3) xor a(4) xor a(5) xor a(1) xor a(7);
end cascade1_arch;

architecture cascade2_arch of gaire_reduced_xor is
	signal p: std_logic_vector(7 downto 0);
begin
	p(0) <= a(0);
	p(1) <= p(0) xor a(1);
	p(2) <= p(2) xor a(2);
	p(3) <= p(2) xor a(3);
	p(4) <= p(3) xor a(4);
	p(5) <= p(4) xor a(5);
	p(6) <= p(5) xor a(6);
	p(7) <= p(6) xor a(7);
	y <= p(7);
end cascade2_arch;

architecture cascade_compact_arch of gaire_reduced_xor is
	constant WIDTH: integer :=8;
	signal p: std_logic_vector(WIDTH-1 downto 0);
begin
	p <= (p(WIDTH-2 downto 0) & '0') xor a;
	y <= p(WIDTH-1);
end cascade_compact_arch; 

architecture tree_arch of gaire_reduced_xor is
begin
	y <= ((a(7) xor a(6)) xor (a(5) xor a(4))) xor ((a(3) xor a(2)) xor (a(1) xor a(0)));
end tree_arch;

